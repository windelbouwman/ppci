../../axi/axi_spi_master/spi_master_clkgen.sv